// $Id: $
// File name:   flex_pts_sr.sv
// Created:     9/13/2015
// Author:      Kyle Rakos
// Lab Section: 337-01
// Version:     1.0  Initial Design Entry
// Description: Flexible parallel to serial shift register
