// $Id: $
// File name:   controller.sv
// Created:     9/28/2015
// Author:      Kyle Rakos
// Lab Section: 337-01
// Version:     1.0  Initial Design Entry
// Description: regulates the controls the operation sequence of the entire system
